module top_module(
    input clk,
    input areset,    // Asynchronous reset to OFF
    input j,
    input k,
    output out); //  

    parameter OFF=0, ON=1; 
    reg state, next_state;

    always @(*) begin
        case(state)
            OFF:begin
                if(j == 1'b1) next_state = ON;
                else next_state = state;
                out = 1'b0;
            end
            ON:begin
                if(k == 1'b1) next_state = OFF;
                else next_state = state;
                out = 1'b1;
            end
        endcase
    end

    always @(posedge clk, posedge areset) begin
        if(areset)begin
           state <= OFF;
        end
        else state <= next_state;
    end
endmodule